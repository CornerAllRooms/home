data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABLAAAAKiCAIAAABJjbIyAAAgAElEQVR4nOzdd3zV9b348c/JIkxBhIIMBRRFEUTAvVCpguM6KlZ/rWIdtbaO2tvbcVvb21Zva3u1lWq1OGrR1gkoIlZEcSIioCIOVIQAMpQ9Qkhyzu+P03tumgQkkJMT8nk+/0q+5zveiT4eebz4rkQqlQoAAADEJy/XAwAAAJAbghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSghAAACBSBbkeAABypHJLKFsdQl5ovkdIJHI9DQDkgCAEIDJr54c5d4aSZ8KquSFZHkIIRW1Ch0PCPl8JfS4MRa1zPR8ANJxEKpXK9QwA0CC2bAgv/3t4588hbOVvX9Fu4ejfhr6XNexYAJAzghCAOKz5KIw/Oayb/8Vr9jo7nPy3UNAs+zMBQI4JQgAisHpeGDskbPx0e9ffa1g4dZwmBKDJ85RRAJq6utZgCGHhpDDxrFBRlrWZAKBREIQANGk7UINpmhCACAhCAJquHa7BNE0IQFPnHkIAGrfyTWHBxDD/8bD6/bBxaShsFVp0Cp0OD91PCnseEwqKt7rhmg/DY8fveA1mfOH9hBuXhpLJYfHz4bM3w+aVIVUZWu8VOgwI+54buhwbEv7tFYDGSxAC0FglK8PbfwzTfxHKVtW+Qn5x6HxU6D40dB8aOgz4l5fL11cNptVswvKNYckLoWRyKJkcVs3d6oa7HxCOuTnsdXL9jAEA9U0QAtAola0NE88Oi5/b3vWL9wjdTgjdhobuQ0NyS33WYNpew8LwR8OquaFkcih5JiydFpJbtnfbQT8OR95Qn8MAQD0RhAA0Pls2hEeOCivf3sHN84rqUGsNs9uDrgxDbqvXaQCgHrixAYDGZ8olO16DIWSlBndyt3NuD+/+pd4mAYB6IggBaGQWPB0+fDjXQ2TBi98NZetyPQQA/AtBCEAjM+OXuZ4gO7asCW+NyvUQAPAvBCEAjcnaT8LSV3M9RNZ8cH+uJwCAfyEIAWhMFj6d6wmyafX7YX1JrocAgP8jCAFoTEom53qCLGvyPyAAuxRBCECjkawMi5/P9RBZJggBaEwEIQCNxoo3wpY1uR4iyxY/F7wBGIBGQxAC0GjEcPas9LPw2Zu5HgIA/kkQAtBoxBCEIYRFcfyYAOwKBCEAjcOWDWHZtFwP0SAi6V4AdgWCEIDGYckLIVme6yEaxKcvh4rNuR4CAEIQhAA0FvGcN6vcHD59OddDAEAIghCA3EulworZYcGTuZ6jAc29K6xbkOshACAkUh5+DUBOrF8cFk0OJZPDomdD6We5niYXdtsndB8aug8NXU8IzXbL9TQAxEgQAtCAtqwPi6f+swNXv5/raRqNRH740uDQbWjoPjR0OjzkF+Z6IABiIQgByL7Nq8Pcu8InE8LSaSFVketpGrfCVqHrkLDviND7qyGvINfTANDECUIAsilZGd64Mcz6XdiyLtej7Gp26xWOuTn0PCPXcwDQlAlCALKmdGV46ithydRcz7ErG/jDcOSNIZHI9RwANE2CEIDsqCgNY08Iy17L9Ry7vsH/GY74Va6HAKBp8toJALLj+W+rwfox44bw8eO5HgKApkkQApAFy6aH9+7N9RBNyEvfDRVluR4CgCZIEAKQBbNvyfUETcu6T8JHj+R6CACaIEEIQH0r3xg+mZDrIZqceQ/megIAmiBBCEB9++zNULEp10M0OUun5XoCAJogQQhAfVv3Sa4naIrKVoWyNbkeAoCmRhACUN8qPf4kOyrLcz0BAE2NIASgvhXvnusJmqhmbXM9AQBNjSAEoL617Z3rCZqiNj1DfmGuhwCgqRGEANS33Q8IzTvmeohcaL132G2fULxHVnbedUhWdgtA3ApyPQAATU4iEbqdGOb9PddzNJS8ojDgurDfBWGPg/655PM54Y3/Dh8+HFKV9XaU7ifV264A4H8lUqlUrmcAoMl5997w7DdyPUSDaN4xnPZ46Hx4LR8teDpMPCtUbq6PwyTCpctDiw71sSsA+D8uGQUgC7oNzfUEDaJt7zBiWu01GELY+5Qw5Pb6OVCHg9UgANkgCAHIgtZdQ7v9cz1ElnU+Mpz7atit57bWOeDi0GabK2ynSAIbgAYnCAHIju5NumF6nR3OmhKat//iNXt/tR4O5wZCALJDEAKQHU34pFb/q8PwR0JB8XatvOfRO3u4/OKw5zE7uxMAqI2njAKQHV2PD4mCkKrI9Rz1KxGO/m045Ht12GLnHzS659HbG58AUEfOEAKQHUWtQ6etPG1lF5XfLJzy97rVYAhh7fydPW7TvvgWgJwShABkTbcTcz1B/WnWLpz5TOh9Xt22SqXCO3fu7KG9kh6ArBGEAGTHuoXhvftyPUQ9ab1XOPeV0OXYOm/40aNh1bs7e/Tp/xUqynZ2JwBQGy+mByAL1i0Mjx0f1i/I9Rz1ocOAcMbE0LJznTdcPiOM+3LYsqYeZtj71DD8sVDQrB52BQBVOEMIQH1rSjXY/eRwzos7UoMLngqPDamfGgwhLJgYnjrHeUIA6p0gBKBeNaUa7HNxOOPJUNSqzhu+MzpMOCNUbKzPYTQhAFkgCAGoP02pBg/9WRh6T8ir+/uZpv00PHd5PbxtoiZNCEB9cw8hAPWkydRgoiCccGc48Bt13rCyPEy5LLyf5UfpuJ8QgPojCAGoD02mBgtbhWGPhL1PqfOGW9aHieeERZOzMFMNmhCAeiIIAdhpG5eGR44O63b6Dew516JTOGNi6HhInTfc8Gl4Ynj4/K0szLQVPc8Mpz4WEm79AGCn+EMCwE6bPLIp1GC7/cOI13akBlfODQ8f3qA1GEKYPz7M/n2DHhGApsgZQgB2zvv3h2e+3hAHShSEPfqFitKweVUoXV7PO9/zmHDa46G4XZ03XDw1PHlWvb1eok7ym4cLPwitu+Xg0AA0FXV/eBoAVDX75qwfolW3cOj1oddZoXn7fy5Z9Fx447/DomfrZ//7nBu+PGZHbsn74O9h8siQ3FI/Y9RVZWmYc0c48obcHB2AJsEZQgB2wsp3wgMHZfcQHQeHf3sqNN+jlo/e+E149Yc7u/+DvxuO+Z+QSNR5w5k3hVd+GEJO/4y26hq+sSiXAwCwi3MPIQA7Yelr2d1/UZvwb5Nqr8EQwqAfhIE7E4R54djfh2NvrnMNppJh6nfCKz/IcQ2GEDYsDhuX5ngGAHZlghCAnbD6/ezuv/9V/3eZaK2OvDHsv0N3MOYXh+EPh4OvqfOGFaVh4jnh7dt25KDZsCrL/wkAaNLcQwjATkhWZHf//a/6ghUSiXDi3WHjsrq9ALC4fTjt8bDnUXWep/TzMOH0sCzL50XrJJXl/wQANGnOEAKwEwpbZHPnrUOLL33xavmF4dTHwh4Hb+9u2/QI576yIzW45uPw8JGNqwZDCAUtcz0BALswQQjATmifzSfK5BVu75pFrcO/PRVa7/3Fa3YcFEZMC+32q/Mwy14PjxwR1n5Y5w2zKxH2yPJDfQBo0gQhADthz6NCqPvzObdT2aqw5uPtXbll5/Bvk0Kz3be1zl7DwzlTt+usYzXzJ4SxQ0LpZ3XeMNs6HByKWud6CAB2YYIQgJ3QunvoPjSL+5/3YB1W3n3/cPqEkF9c+6cHXhZOfyIU1v0Cyzl3hIlnhYpNdd6wARx4Wa4nAGDXJggB2DmD/zOLJwnn/CmUfl6H9fc8Mpzy91r+uh3+y3Din0Neft2OnkqFV34Unv9WSFXWbcOG0Xqv0OfCXA8BwK5NEAKwc7ocGw66Ils737gkPPWVUFFWh016nRmOH/V/3+YVhqH3hUN/UudDV24Jz3w9zPx1nTdsMCeO3pETngBQhSAEYKcdc0voekK2dr7khTD5opCqyyvg+135zxfWF7UJZzy1I6fRytaGx4eFDx6o84YN5ujfZfdiXQDikEjV6U8sANSqfFN4YnhY8kK29j/gunDM/9Rtk5f+Pez/9dChf52PtX5xeGJ4WDmnzhs2mCN/HQb9INdDANAUCEIA6km2m/CYm8OA72Zr5xmfzwmPDwsbl2T9QDtMDQJQfwQhAPUnu02YCKf8PfQ+Lzs7DyGEsOi5MPHssGVtFg+xk9QgAPVKEAJQr7LahPnNwr/9I3Q9Lis7f//+8Ow3QrI8KzuvF2oQgPrmoTIA1KvCFuGMiaFLdpqtsiw8eWZY+U7973nGjeGZC9UgALFxhhCALCjfGJ44NVvnCVt1DedOC6271s/ekpVh6nfCO3fUz96yRA0CkB2CEIDsKN8YHh8WPn0pKzvfvW849+XQbLed3U/5pvD0V8MnE+pjpqw54oYw+Me5HgKApsklowBkR2HL0OGQbO181TvhyTPr9sL6mjatCI8d39hrMITQ6bBcTwBAkyUIAciaRZOzuPMlU+v8wvqq1nwYHjkyrJhRrzNlR8mzuZ4AgCZLEAKQHRuWhFXvZvcQHz4UXvrejmy4dFp4+Miw9uP6Hig7strVAMRNEAKQHYsa5LzWm7eEWTfXbZOPx4exJ4bNn2dnoCxYMTuUrsz1EAA0TYIQgOwoaajzWi//e5j30Pau/NYfw8RzQmVpNgeqd8mwaEquZwCgaRKEAGRBKtWAd76lwuSLwuKpX7RWKrz8/fDCVSEkG2Ko+uWqUQCyQxACkAUr54TS5Q13uPQL6z+fs/UVtoSnLwizftdwI9WvBjvdCkBkBCEAWdDwAbNlbRh3Ylg2vZaPNq0I44aGDx9s6JHq0fqFYc2HuR4CgCaoINcDANAUNcwTZaop/Sw8fETY5yuh7+Vh9wNCQXFY+3F4f0x4/4FQtioH89Svksmh7b65HgKApiaR2uE3OAFArSq3hDvbhYpNuZ6jael5ZjhtXK6HAKCpcckoAPVtxSw1WP8+fSnXEwDQBAlCAOrbuvm5nqAp2rwylMtsAOqZIASAXUTZmlxPAEBTIwgBqG+J/FxP0EQVt8v1BAA0NYIQgPrW/qBcT9AUtegcCprneggAmhpBCEB9a39AaLlnrodocroPzfUEADRBghCALOh1Vq4naHJ6fzXXEwDQBAlCALLg0OtDUZtcD9GEdBwY9jol10MA0AQJQgCyoEXHcOj1uR6iqcgvDifcGRKJXM8BQBMkCAHIjgHXhf0vzPUQTUAifPmvoePAXI8BQNMkCAHIjkQiDL03HHxtCE5t7aii3cKpY8O+5+Z6DgCarEQqlcr1DAA0acteDy9cHZZPz/Ucu5a80Pur4Yhfht165noSAJoyQQhA9qVSYdlrYf4ToeSZ8NnsEPzp2Yr84rDn0aH7l0Ovs0PbXrmeBoCmTxAC0LBKPw+LpoSSyaFkcthQkutpGoNE6HBw6HZS6D407HlMKCjO9TwAREQQApA7q+eFkslh0eSweGrYsjbX0zSsVt1C96Gh+9DQ9cTQokOupwEgUoIQgEYgWRkePiKsmJHrORrKIf8Rjv5NrocAAE8ZBaAxyMuP68XrPU7L9QQAEIIgBKCx6D401xM0lMJWodPhuR4CAEIQhAA0Fp0OD4Wtcj1Eg+hyfMgvzPUQABCCIASgscgvDF2Oy/UQDSKec6EANHqCEIBGI5JSiuTHBGBXIAgBaDS6RVBKLbuE3fvkeggA+CdBCECj0f6A0LJLrofIMqcHAWhMBCEAjUm3k3I9QZYJQgAaE0EIQGPSxHsp0fSLF4BdiiAEoDHZ6+SQyM/1EFnTYUBo0THXQwDA/xGEADQmzfcIPU7P9RBZc9A3cz0BAPwLQQhAI3P0TSGvKNdDZEHrvUKfkbkeAgD+hSAEoJFpu2845Hu5HqK+JQrCyfeH/KYYugDsygQhAI3PEb8K+563g9u26RHaH1Sv0/yvzkeFwtY7tGVeGHJ72PPoep4HAHZaIpVK5XoGAKghlQwvXhfeGhVC8otXLmobup0Qug8N3YaGtr1C+aYw4fSw+Ln6nOew/wqHXR+SFWHZ9FAyOSyaHJa9HlIVX7xhYevw5b+GXmfW5zAAUE8EIQCN2PI3wrSfhJLJtWRhXmHodEToPjR0Hxo6Dgp5//ps0vptwnQNVlO2Lix+PiyaHEomhzXzatkqvzjsd0E4/BehVZf6GQMA6psgBKDR27g0fDIhrJ4XNn4aCluFFl8KnY8Iex4bilpta6v6asJaa7Ca9SVh0XPhs9lh88qQrAht9g579A89TgtFO3aJKQA0EEEIQNO18024PTUIALssD5UBoOkqbBFOnxC6nrCDm6tBAJo6QQhAk7bDTagGAYiAIASgqduBJlSDAMTBPYQAxKFic5h8cfjwwS9YLb9ZOOq34eCrGmQmAMgxQQhATD58NLz6w7D249o/7XpiOO7W0P6Ahp0JAHJGEAIQmVQqLHo2LPxH+Gx22LQsJPLDbr1Cx0PCviNCu/1yPRwANChBCAAAECkPlQEAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIhUQa4HAIDozJ49+29/+9usWbNWrlzZokWL008//Qc/+EFe3o78K+3MmTMXLVqUSqUSiUT//v179OhR79MC0IQJQgC+WGVl5XvvvTd37tw1a9YUFxf37NnzkEMOadmyZa7n2vVUVFT89re/veGGGzZu3JhekkgkunTpkkqldmBvlZWVt95665gxY1KpVH5+/i233HLVVVfV67wANHEuGQVgWzZs2HDzzTf36dOnX79+X/3qV6+44oqRI0ced9xx3bp1u+qqqz799NNcD7iLmTJlyk033ZSpwSxJJpO//OUvi4qKCgoKioqK/ud//ierhwNg1+UMIQBbNX/+/EsuueTFF19MJpNVl6dSqdWrV992222vvPLK/ffff8ABB+Rqwl1LMpl88skn165dG0JIJBJ9+/a94YYbBg8enJeXl5+fX48HysvLKygoqKysTP+HKyjw5x6A2vkLAUDt1qxZc/XVV7/wwgvpqxlbtmx56KGHdu7cef78+bNmzdqyZUsqlXrzzTevu+66v//97+3atcv1vLuALVu2fPLJJ+nfZ0FBwTXXXHP66adn6VhFRUWJRCLzdZaOAsCuziWjANRuypQpzz//fLpe9txzz/Hjxz/33HMPPPDAK6+88sADD+yxxx4hhFQq9cILLzz55JO5HnbXUF5evnnz5vTXhYWFu+++e/aOVVhYmPlaEAKwNc4QAlCLZDL52muvpeslkUgceeSRxx9/fPqjvLy8s84667XXXrvllluSyWRZWdmTTz553nnnFRUVzZgx45VXXsk88XLIkCFV97l+/fqxY8euWrUqhNCyZcuzzjqrQ4cOVVdYvXr1uHHjpkyZsnDhwrKysg4dOgwcOHDEiBEHHXRQrUNWVFQ8//zzEyZMmDt37tq1a1u3bt27d+/TTjvt5JNP3loCzZs377HHHps+ffrSpUuTyWS3bt2OO+648847r1OnTjVXXrNmzdixY6dMmbJgwYKysrJ27doNGDBgxIgRgwYNqrnyBx988NBDD82YMWPZsmWJRKJr167HHHPM+eefn9nzvHnzZsyY8dlnn6W/raysfOONNyoqKhKJxIABA7p16/bEE08sWrQohFBUVDRs2LCePXtW3f9HH300adKkioqKEMLee+991lln1foDZmR+A4lEomocAsC/SAFADRUVFZdcckn6msNEInH22WeXlZVVXeHpp5/u1atX586dO3fuPHTo0OXLl6dSqRtvvDH97oREIvGtb32rsrKy6iYLFizo3bt3+q9Pp06dZs+eXfVw999//9577525yjGjuLj429/+9sqVK6tN+NZbbw0ZMqTmrXd5eXlHH3101Z2nrVu37j/+4z/atGlTbf30Qz7HjBlTbdqJEyf27t275jwtWrT4/ve/v2HDhsyapaWlP//5z2vdc7du3R599NH0ajfddFOtL5bIz8//wx/+sGbNmkw/t2zZ8vHHH682/8MPP1xcXJxe4ZRTTsn83i688ML0kPn5+bfeemtm/bvvvjv9yyksLHzggQe+4L83ALFyhhCAWiQSiXbt2iUSifRfi2nTpr366quZk4QhhJNPPvmjjz6ql2NVVFTcdNNNv/rVr0pLS2t+unnz5j/96U9Lly69++6727Ztm174wgsvXHTRRSUlJakab2tIJpOvvPLKOeec89BDD2VO5a1cufKKK64YN25cZWVltfVTqdSSJUu+/e1vV1ZWXnTRRemF06dPv/zyy5csWRJCyMvLa9++fWFh4fLlyysrKzdt2vT73/++efPm119/fX5+fjKZHDVq1I033rhly5YQQmFhYadOndavX7927dpUKrVo0aIrr7yyXbt2J5xwQr38rrZfYWFhXl5eZWVl+gEzDXx0AHYV7iEEoBZ5eXmDBw9u1qxZ+ttly5ade+65P/zhD999991qTxzdeU888cRvfvObdA22adPmZz/7WUlJycqVK+++++4uXbqEEJLJ5IQJE+666670+gsXLrz22mvTNZifn3/WWWe98cYbGzZsePHFF48//vh0xH7yySfXX399+nmeFRUVv/71r9M1mEgkBg0aNHHixHXr1n388cfXXntt+rTbunXrfvGLX7zzzjvpw40ZMyb9Ro28vLxLL730k08+KSkpGT16dPo0YHl5+b333vvuu++mfzP3339/ugbbtGlz3333LViw4JNPPrn44ovT5wM/++yzUaNGbdq0afjw4X/6058OPPDA9E/RrFmz7373u/fcc89dd901dOjQ+v2VhipPFhWEAGyDIASgdieddNKxxx6bvhwxlUp9/vnnv/nNb/r167fffvtdcskl48eP37Rp084fZfXq1aNGjVq/fn0IobCw8Pvf//7111/frVu33Xff/Rvf+MZ///d/t2jRIoRQXl7+0EMPLV++PJlM/vWvf50zZ04qlUokEscff/zo0aMHDhzYsmXLY4455o477khflZpKpV599dXXX389hDBr1qwHHnggfW6wZ8+e99577/Dhw1u3bt2zZ89f//rX559/fvpnXLBgwZgxY5LJ5KZNmz744IP0ucfCwsITTjihZcuW+fn555133nHHHZdeedmyZTNmzAghLFmyZNmyZemfpVOnTkcccUReXl7btm2vueaazp07pyeZNWtWSUnJgQceeP7553fs2DG9ckFBwXHHHXfxxRePHDmyT58+O/+brKagoCB9yaggBGAbBCEAtdt9993vuOOOYcOGVb1Pr7Ky8qOPPrrnnnvOPvvsfv36jR49uqysbGeO8tZbb7355pvp+tp7773PP//8qjfanUwao7MAACAASURBVHDCCfvss0/664ULFy5YsGD16tWTJk1K111RUdHIkSPbt2+fWX+fffY54YQT0s22fv36mTNnJpPJiRMnLl++PISQSCROPfXUqm9NbNas2bnnntu6desQQjKZfP755z///POqbwXcsmXL+PHj16xZE0Jo0aLF3//+988++2zFihVLly694IILwv9emZleefHixU8//XR6tr59+77zzjsrVqxYsWLF7Nmz99133535Le2AgoKC9GCCEIBt8BcCgK3ae++9x40bN27cuNtuu+21114rLy/PfJRKpT7++OMrr7xy+vTpt9xyS7qpdsCcOXPSpwcTicQ+++yTPquW0blz53HjxqVXyM/P33vvvT/++OOFCxemP919992rPYA0Pz//v/7rv6644or0+cMOHTps3rz5jTfeSAdnfn5+UVHRxIkTq26yfPny4uLidevWhf893de3b9+BAwdOnjw5mUymUqmHHnpo5syZI0aMOO200wYNGtSyZcuqm3fp0qVHjx7pZ+ps2rTp6quvfuihh0aMGHHKKaf06NFjx34n9aJqEHrKKABbIwgB2JaioqLzzjvvvPPOmzdv3qRJk5577rkXX3wx/cSUEEJFRcVf//rXHj16/OhHP6r1EZrblkwmFy9enHkwTPv27TN3Labl5eVVe/vCZ599lrlUtVWrVrvttlu1fXbo0KHq2yxWrFjx2WefZab93e9+97vf/W5r85SWlq5ZsyYvL+8b3/jG008/nXlU6YcffnjDDTfceOONXbp0Ofvss6+88sr99tsvc7hrr732m9/8ZvosYnl5+dSpU6dOnVpYWNivX7+LLrrowgsvrDlkA8gEoddOALANLhkFYLv07t37mmuuefzxx+fPn/+rX/0q81L18vLyBx98MP1Azm2r+UTQEMLmzZszy7fnysaysrLMk0ITiUTN10JUU1lZmX5333ZKD9OrV6+xY8deeOGF6TsYMx8tXrz41ltvPfLII//85z9nxhgxYsQjjzxy2GGHVb22try8fObMmddcc82QIUNmzpy5/QNsTfp05favn7mWteoVsABQjTOEANRNu3btfvzjH7dv3/7aa69Nv7l+8eLFH330Ubdu3aquVjPDtmzZkl6/qhYtWqSfCxpCWL9+/Rc2T/PmzTN5s3nz5i+8g7GgoCBz1rFFixZXXXVV5uReTcXFxZk7DPfaa6+//OUv119//fjx45955plp06Zlxlu1atUPf/jD7t27n3LKKemVTzrppCFDhkybNu2JJ56YMmXKnDlz0pfXplKpN99889vf/vb48eMzb6j/QqlUqubrMUpLS2su3PYPnnk/oTOEAGyNIASgFnfddddPf/rT9HsajjrqqPvuu6/aXYJDhgz50pe+lL6dr7y8PPOY0MwK69atq1Z3n376aXq1jLy8vO7du+fl5aVPfy1ZsmTt2rVVHxKzefPm5557buXKlSGEZs2aHX/88R07dmzZsmX6+sx169YtWbIk87L7tJkzZ7733nvpewj79+/fu3fvjh07ppuzvLx8//33HzlyZLUftqKiIv0ujfz8/Gon03r27Hndddddd911q1atGj169O9+97vPP/88hLBmzZpHH3106NChmfXz8/OPPvroo48+OoQwd+7cX//61w899FB5eXkqlXr77bfTr0bcxi+86qHLy8s3btxY9dNkMvnxxx/X6YUfBx100F/+8peysrLi4uJtNDAAkROEANSiW7dumzZtSj9q5fnnn3/55ZeHDRtWdYXS0tLMM2aKiorSt8mlT/eF/33b+9q1azNXliaTyalTp6Z3WFXfvn3btGmzatWqEMK8efPmzp177LHHZj595513Lr300qVLl4YQevXq9Y9//KNLly49e/ZMX6G6fv36qVOnHnfccZnbF9evX/+f//mfzzzzTCqVKioquvvuuw866KD0iwfT144+99xzF1xwQVFRUeYQEyZMuOCCCzZs2JBIJI499tjx48e/8cYbf/jDH9IxfOihh/7oRz8qKirafffdf/CDH+Tn5//oRz+qqKhIv3R+48aNo0aNevXVV9NvRLziiitOPfXUEMKBBx54++23r1ixYvLkyalUasuWLSUlJdv+hVc9k1lZWfnhhx8mk8nMz7VmzZoXXnihTpeMtm/ffvjw4atWrWrfvr1LRgHYGvcQAlCLQw455IADDkjX3dq1a6+99trnnnsu8+nKlSt/+9vfZt6/t/fee6dP03Xs2DFzkvDtt99+5plnMptMmzbt3nvvrXnRY79+/QYOHJg+0OrVq2+66ab0+cAQwvr163//+9+nj5JIJI4++uhu3bq1a9futNNOS99tWFlZee+9906bNi29fjKZfPDBB19++eV0OPXo0eOII44IIZxyyilf+tKXQgipVOrJJ5+cMGFC5ugrVqy47bbb0qfj8vPzhw0b1rZt22bNmk2bNm3SpElPPfXUn//851mzZmXW32233dKjJhKJZs2aFRQUVFRU/OMf/5g0adLEiRNHjRq1evXq9JpFRUWZ55EmEoni4uJt/8ILCws7deqUyelx48bNnz8//VFlZeVdd931+uuv1xqEmdhLpVLpE6dpL7300oEHHti5c+f+/ftPnz5920cHIFrOEAJQi/TDMy+//PL0lZ/z5s0bNmzYgAEDevfuvWHDhunTpy9dujTdJ8XFxZdddln6dREHH3xw9+7d582bF0JYt27d5ZdfPn78+D59+ixatGj8+PGVlZWtWrXasGFD1QPttttu11577cyZM1etWpVKpSZNmjRkyJAzzjgjPz9/0qRJM2fOTB+lS5cuV155ZfrM3te+9rVx48ZNnz49/ZSXM88885xzztlrr71mzZo1ceLE0tLSEEJRUdFll12WfvHDIYccMnLkyJtuuqmiomL16tUjR4585JFH+vfvv2bNmieeeCL9DvpEIjFgwICvfe1r6Z/iqKOOmjBhQiqVWrp06f/7f//vW9/6Vp8+febNm3frrbem743Mz88/8sgjW7RoccYZZ9x9992LFi1KpVLPPvvsueeeO3LkyDZt2jzzzDPpE5UhhPbt2w8YMGDbv/D8/Pzjjz/+gQceSD9l55133hk6dOjpp5/erl27119//bnnnmvXrt3KlSur3ZmZSCSaN2+e/jqZTN5yyy2zZ8/+6U9/2qdPn5tvvvnDDz9MpVLvvvvuLbfc8uCDD9bH/xcANDkpAKhNRUXFH//4x7Zt227jj0jLli1//vOfpxsmlUpVVlbedtttVZ/MmVFUVPT9738/c79fp06dMi91qKysHD16dLt27bZ2lI4dOz788MNVZ5s9e3b//v239ojRwsLCa665ZuPGjZn1161bd8UVV2zt2SqJROKAAw6YMWNGZv0333yzT58+W9t/IpEYOnRoOokrKyvvuOOONm3abG34oqKin//85+mbCdetWzdkyJDMr278+PFVf6g1a9aMGDGi1rd3dO3a9ac//WnmNOMpp5yS2er222+v+nO1adPmqaeeWrdu3YknnpiZdvjw4fX8PwcATYUgBGBbZs2adcEFF2QulcwoLi4+9dRTX3zxxWrrV1RU3HfffT179sysn0gk2rRpc/XVV8+ZM6fWIEx7+eWXTz755GrN1rJly/POO2/OnDk1B1uyZMnVV1/drl27qoPl5+cPHjz4kUceSd/mV1VZWdmYMWP69etXtbgSiUTHjh2vu+66dN1VtWDBgssvv7xt27ZV959IJPbcc8/rr79+5cqVVVeeMmXKkCFDqg2fn58/cODAzKNlUl8UhKlUauXKlddee22bNm2q/vZ69Ohx3333Pfjgg7UG4cqVKy+++OLM/YfpIEylUrfffnu6zFu1anXPPfds+78yANH655O+AWAbNm7cOHv27I8//njdunXFxcVdu3YdOHBgx44dt7b+5s2bZ8yY8cEHH5SXl3ft2vXwww+v+rL4bViyZMmMGTOWL1+efgDpoEGDqj50tNbBpk+fvmDBgi1btrRv3/6QQw7p0aNHrSfZ0pLJ5Pvvv//222+vXr26uLh43333HTBgQOZmv5rWrl07e/bs+fPnl5aWtmrVar/99hswYECmvqopKSmZPXv2smXLksnkHnvs0b9//3322Wcbw2zNihUrpk2btmTJkqKioj59+gwaNGhrR8xYvnz5woULU6lUmzZtevToUVxcnEwmX3/99bfffnvAgAEDBw7cgTEAiIEgBAAAiJR/LwQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIiUIAQAAIhUQa4HAICGUFlZ+e67786YMeONN96YOXPmypUrS0tLN2/enEgkmjdv3rx5865duw4aNGjw4MGDBg3q0aNHrucFgIaQSKVSuZ4BALJl4cKFo0ePnjp16uzZszdt2rSdW+2xxx6DBg0aNmzYyJEj27Rpk9UJASCHBCEATdOUKVNGjRo1YcKEZDK5wztp1arV17/+9e985zsHHHBAPc4GAI2EIASgSSkrK7v77rv/+Mc/vvfee/W42xNOOOGaa64544wz6nGfAJBzghCApmPWrFkXXnjh3Llzs7T/008//c9//nOnTp2ytH8AaGCeMgpAU1BeXv6zn/3ssMMOy14NhhAmTJjQt2/fBx98MHuHAICG5AwhALu8OXPmXHTRRbNnz/7CNVu3bj1w4MBBgwYdeOCBLVu2LC4uTiaTmzdvXrNmzZtvvjljxoy33367vLz8C/dz7rnn3n777XvssUd9jA8AOSMIAdi1jR079vzzz9+yZcs21jnssMMuvfTSo446ar/99svL29bVMWVlZW+//faUKVPuvPPOBQsWbGPNPffcc8qUKfvvv/+OjQ0AjYEgBGAXNnbs2K9+9atbO6fXrFmzESNGXHXVVYMHD67rnpPJ5IQJE/74xz8+++yzW1unU6dOzz//vCYEYNclCAHYVW27Bi+99NIbb7yxQ4cOO3mUuXPnfutb33rppZdq/VQTArBLE4QA7JK2UYNdunQZPXr0sGHD6utYyWTyD3/4w49//OPNmzfX/FQTArDrEoQA7HqmTJkybNiwWmvwa1/72qhRo9q2bVvvB/3ggw8uuuii6dOn1/yoU6dOM2fO3HPPPev9oACQVYIQgF3M2rVr+/btu3jx4pof3XDDDT/+8Y+zd+jy8vKvfOUrTzzxRM2Phg8fPnHixOwdGgCywXsIAdjFXHPNNTmpwRBCYWHho48+esYZZ9T86Kmnnrr77ruzenQAqHfOEAKwK5kwYUKtPdYANZixtfOEbdq0mTNnTvfu3RtmDADYeYIQgF3GypUr+/btu2zZsmrL//3f//23v/1tQ05SXl5+0kknvfjii9WWn3jiiZMnT04kEg05DADsMJeMArDL+OEPf1izBvv163fDDTc08CSFhYV/+ctfWrVqVW35lClTxowZ08DDAMAOc4YQgF3D559/3q1bt2ovfigsLJwxY0b//v1zMtKdd955xRVXVFt48MEHz549OyfzAEBdOUMIwK5h9OjRNV8DeP311+eqBkMI3/zmN08++eRqC998882XX345J/MAQF05QwjALqCysrJHjx6LFi2qurB3795z584tKCjI1VQhhJKSkl69elVUVFRdOGLEiIceeihXIwHA9nOGEIBdwPjx46vVYAjhO9/5Tm5rMITQvXv3s846q9rCsWPHLlmyJCfzAECdOEMIwC5gyJAhU6dOrbqkdevWS5Ysad269Ta2qqiomDZt2oIFC9avX59MJlu0aLHPPvsMGDBg21t9/vnnr7766ltvvbV+/fri4uIDDjjgiCOO2Guvvba2/ksvvXTsscdWW/iTn/zkl7/85Rf/YACQU4IQgMZu7dq17dq1q/YH6zvf+c6oUaO2tsmUKVPuueeeSZMmrV69utpHiUTioIMOGjduXM+ePat9NH/+/Ouvv/6RRx7ZsmVLtU2GDh36i1/84rDDDqv1cAcffPBbb71VdUm/fv2qLQGARkgQAtDYTZky5aSTTqq28L333tt///1rrrxs2bJLLrnkqaee2sYOCwsLV69e3bJly6oLH3vssYsvvnj9+vVb26qgoOA3v/nNddddV/Oju+6667LLLqu6JD8/f/369c2bN9/GGACQc+4hBKCxmzFjRrUle+21V601OG/evCOOOGLbNRhCOPTQQ6vV4NSpU88///yqNdi2bdtevXpVvbi0oqLie9/73t/+9reaO6z5rNHKykovnwCg8ROEADR2NYNw0KBBNVfbuHHjGWecsWDBgsySrl27XnfddS+99NLChQtLSkrmzJkzZsyYK6+88itf+UrVDRcuXHjOOeeUl5env91tt91uvvnmFStWfPTRRytWrPjlL3/ZokWLzMqXXnrpnDlzqh26W7duX/rSl75wbABobHL8cDYA+EJvvPFGtSWDBw+uudpPfvKTDz74IPPtl7/85bFjx1Y9E9itW7e+fft+7Wtfq7bhnXfeuWrVqsy3Y8aMOf3009NfFxcX/+QnP+nevftFF12UXlJaWnrHHXfcdttt1XYyaNCgiRMnVl0iCAFo/JwhBKBRW7FiRUlJSbWFNYNw7dq1d911V+bbY4455sknn6x2XWitUqlU1atAzz///EwNZlx44YVVLwp99NFHKysrv3AkQQhA4ycIAWjUql4CmnHIIYdUW/L4449v2LAh8+33vve9wsLC7dn/yy+/vHDhwsy35557bq2rnX/++ZmvV6xYUe0dGLWOVHW3ANA4uWQUgEattLS02pK8vLy2bdtWW1j1stJOnTqddtppmW/Ly8s//PDDausXFBT07t07hPCPf/yj6p6PP/74Wseo9pjT11577cQTT6y6pH379tU2KSsrSyaTeXn+7RWAxksQAtCo1QzCWt/l8P7772e+7tWrV35+fubbkpKSAw88sNr6HTt2XL58eQih6t2D7dq1a9euXa1jdOnSpbCwMPPgmZpvp6h1qtLS0u25bBUAcsU/WwLQqNW8W69q7GVs3rw583VRUdH277+srCzz9bavMi0o+L9/Ra35Ft9ap6o5PAA0KoIQgEatuLi42pKa5wxDCFXfDLFy5crt33/VM3jr16+vWXppmzdvrtqcbdq02Z6pvJgegEZOEALQqNVsqvLy8oqKimoLO3XqlPl6zpw5n3zySebbbt26zZkzZ86cObW+U7579+6Zrzdu3PjWW2/VOsarr75atRX32muvaits2rSp2pL8/PztfLANAOSKIASgUav1pr6qdwymnXnmmZmvU6nUfffdl/m2qKiob9++ffv27dmzZ81dnXPOOVW/feaZZ2od49lnn818XVhYWPWhNVsbqeaTbwCgsRGEADRqvXv3rno5aFrNV/wNHz68aoDddNNNU6ZM2Z799+jR49BDD818e8stt3z++efV1ikpKan6JvohQ4bUjL2aI9V8EQUANDaCEIBGLT8/v2ZZ1ayvoqKia665JvNtaWnp6aeffuedd9Z8HGhNF1xwQebrZcuWff3rX6/66NHly5d//etfX7duXWbJd7/73Zo7qTlSzVfVA0Bjk9ja3fMA0Ehcd911t9xyS9UlgwcPfv3116utVl5efvjhh8+aNavqwpYtWw4dOrR9+/bl5eVz5syZPXv2/2/v/kJr/v8Ajn9amU5bh4jMn4ii5U8Ni9A04UJSQpbyt0iZFEr5k1rElQsUsciFduF/KCKTQkwJQ7ughCYaF/4czhx9L9S309ns5+s3Zzt7Px6Xr/M5n8/7XK3neZ99Pj/n/z524ucbZ86cmf6s+R49eqxcuXLAgAGvXr06dOhQelVWVFTU1NRkXPrLly/xeDzjnqKnT5+eO3fuH3xeAMgaQQhAZ1dTU5O+iRdFUX5+/ocPH1r+lPTdu3ezZs1Kf0j9r6QHYRRFTU1NEyZMePbsWdvvmjZt2sWLF1ve+PT69evl5eUZw5cvXw4cOPB/rgQAOpCfjALQ2bX87WUymTx+/HjLI/v06XPz5s3du3f36NGj7XNm3Kumd+/edXV18+fP/9Xx3bp127p166VLl1rWYBRFR44cyZj069dPDQLQ+dkhBCAH9O/fv7GxMX0yevTohw8f/ur45ubmGzdunD9//t69e58+fUokEt27d+/Zs+eoUaNKSkpKSkrGjh2bl9fKt6IPHjyorq6+c+dOQ0NDKpWKx+NDhw6tqKhYuHBhnz59Wr3W27dvBw0alEwm04fz588/ceLEH31WAMgeQQhADti+fXtVVVXG8Pr161OnTu2Q9aTbsWPHtm3bMoZXrlyZPn16h6wHAH6fIAQgBzQ2Ng4ePLi5uTl92Bl24b5//z5kyJDXr1+nD4uLi588edJRSwKA3+d/CAHIAUVFRRlPkI+i6MyZM3fu3OmQ9fxr//79GTUYRVFlZWWHLAYA/is7hADkhlu3bk2ePDljOGLEiPv378disQ5ZUkNDQ0lJSSKRSB/G4/HXr18XFhZ2yJIA4D+xQwhAbpg0aVLLJ9Q3NDRs2bKlQ9aTSqWWLl2aUYNRFC1fvlwNApAr7BACkDOuXr06Y8aMjGFeXl5tbW1ZWVmWF7Nr167NmzdnDHv16lVfX19UVJTlxQDAn7FDCEDOmD59+urVqzOGP378qKioaGhoyOZKzp07t3379pbzffv2qUEAcogdQgByyefPn8eMGfP8+fOMeVFRUW1t7YgRI7KwhnPnzi1YsCDjlqdRFM2bN+/kyZNZWAAAtBdBCECOuXHjRnl5+Y8fPzLm2WnCX9Vg37596+vrf/XwegDonPxkFIAcU1ZWtm7dupbzxsbG8vLy27dv/71LHz16tNUajKLo4MGDahCAnCMIAcg9u3fvnj17dst5Y2PjlClTNm3a9O3bt/a94ps3b+bMmbNixYpWa7Cqqmru3Lnte0UAyAI/GQUgJyWTyXnz5l24cKHVV0eOHHns2LFx48a1y7VqamoqKyvfv3/f6qtVVVXbtm1rlwsBQJbZIQQgJ+Xn5586darVfcIoih4/fjxx4sTFixffvXv3jy+RSqXOnj07bdq0RYsWqUEAuiQ7hADksLb3CX8qLS1du3btwoUL8/Pzf/O0TU1N1dXVBw4cePHiRRuHqUEAcp0gBCC3JZPJjRs37t+/v+2/aPF4fNy4caWlpaWlpePHjx8yZEj6q6lU6unTp3V1dXV1dffu3Xvw4EEymWzjbAUFBXv27Fm1alW7fAQA6CiCEICuoLa2dvny5W1v6KUrKCgoKCiIxWKpVCqRSHz69On370NTVlZ29OjRoUOH/uliAaCzEIQAdBEfP37csGHD4cOH/94lYrHYzp07161bl5fnn/AB6AoEIQBdyuXLl9evX//kyZN2P/PMmTP37t37tx98DwDZJAgB6IKuXbu2b9++8+fPp1Kp//NUhYWFS5YsqaysLC4ubpe1AUDnIQgB6LJevHhx4MCB6urqpqamP3j78OHD16xZs2zZsng83u5rA4DOQBAC0MV9//69vr7+5+1D6+rq6uvrm5ubWz2ysLBw7Nix48eP/3kz0mHDhmV5qQCQZYIQgLB8/fr10aNHTU1NiUQikUjk5eXFYrFYLDZgwIDi4mJ3iwEgKIIQAAAgUL4HBQAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAAYweLVQAAAP1JREFUCJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACJQgBAAACNQ/xn2tRJO2KKcAAAAASUVORK5CYII=
